
--------------------------
--addr from pe added as new input
---------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library work;
use work.Pack.all;

entity ControlSignals is
	port (reset: in std_logic;
			IR: in std_logic_vector(15 downto 0);
	      done: in std_logic;
	      addr: in std_logic_vector(2 downto 0);
	      M8_Control_PE: in std_logic;
	      HDU_output_PC: in std_logic;
	      HDU_output_M3: in std_logic;
	      HDU_output_IF_ID: in std_logic;
	      --FDU_output: in std_logic;
	      M2: out std_logic;
	      PC_write: out std_logic;
	      IF_ID_Write: out std_logic;
	      M1: out std_logic;	   
	      M3: out std_logic;
	      M4: out std_logic;
	      M5: out std_logic;
	      M6: out std_logic;
	      M7: out std_logic_vector(1 downto 0);
	      M8: out std_logic;
	      M9: out std_logic_vector(1 downto 0);
	      M10: out std_logic_vector(1 downto 0);
	      --M11: out std_logic_vector(1 downto 0);
	      --M12: out std_logic_vector(1 downto 0);
	      M13: out std_logic_vector(1 downto 0);
	      ALU_OP: out std_logic_vector(1 downto 0);
	      C_en: out std_logic;
	      Z_en: out std_logic;
	      M14: out std_logic;
	      M15: out std_logic;
	      M16: out std_logic_vector(1 downto 0);
	      M17: out std_logic_vector(1 downto 0);
	      M18: out std_logic;
	      M19: out std_logic;
	      M20: out std_logic;
	      Mem_en: out std_logic;
	      Mem_R_W: out std_logic;
	      RF_Write: out std_logic;
	      clk: in std_logic);
end entity;

architecture Behave of ControlSignals is
signal PC_write_tem: std_logic := '1';
signal M2_tem : std_logic := '1';
signal IF_ID_Write_tem : std_logic := '1';
signal M3_tem :std_logic := '1';
signal tm20: std_logic := '0';
begin

    process(IR,done,addr,M8_Control_PE,HDU_output_PC,HDU_output_M3,HDU_output_IF_ID,reset)
		
    begin
         tm20 <= '0';
			M2_tem <= done;
			PC_write_tem <= (done and HDU_output_PC);
			IF_ID_Write_tem <= HDU_output_IF_ID;
			M3_tem <= HDU_output_M3;
		if(reset = '1') then
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '1';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '0';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		else	
		if(IR(15) = '0' and IR(14) = '0' and IR(13) = '0' and IR(12) = '0' and IR(1) = '0' and IR(0) = '0') then ---add
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '1';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '0' and IR(12) = '0' and IR(1) = '1' and IR(0) = '0') then---adc
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '1';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '0' and IR(12) = '0' and IR(1) = '0' and IR(0) = '1') then---adz
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '1';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '0' and IR(12) = '1') then---adi
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '1';
			M9(1) <= '1';
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= '0';
			--M11(1) <= '0';
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '1';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '1' and IR(12) = '0' and IR(1) = '0' and IR(0) = '0') then---ndu
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '1';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '1' and IR(12) = '0' and IR(1) = '1' and IR(0) = '0') then---ndc
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '1';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '1' and IR(12) = '0' and IR(1) = '0' and IR(0) = '1') then---ndz
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '1';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '1' and IR(14) = '1' and IR(13) = '0' and IR(12) = '0') then---beq
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '1';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '1';
			C_en <= '0';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '0';
			M16(0) <= '0'; --depends on alu(zero flag set?)
			M16(1) <= '0'; --depends on alu(zero flag set?)
			M1 <= '1';
		--end if;

		elsif(IR(15) = '1' and IR(14) = '0' and IR(13) = '0' and IR(12) = '1') then---jlr
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7(0) <= '0';
			M7(1) <= '1';
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= '0';
			M10(0) <= '0';
			M10(1) <= '0';
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '0';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '0';
			M17(0) <= '0';
			M17(1) <= '1';
			M18 <= '1';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0'; 
			M16(1) <= '0'; 
			M1 <= '1';
		--end if;

		elsif(IR(15) = '1' and IR(14) = '0' and IR(13) = '0' and IR(12) = '0') then---jal
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			M3_tem <= '0';
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7(0) <= '0';
			M7(1) <= '1';
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= '1';
			M10(0) <= '1';
			M10(1) <= '0';
			--M11(0) <= '0';
			--M11(1) <= '0';
			--M12(0) <= '0';
			--M12(1) <= '0';
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '0';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0'; 
			M16(1) <= '0'; 
			M1 <= '1';
		--end if;

		elsif(IR(15) = '0' and IR(14) = '0' and IR(13) = '1' and IR(12) = '1') then---lhi
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7(0) <= '1';
			M7(1) <= '0';
			M8 <= M8_Control_PE;
			M9(0) <= '1';
			M9(1) <= '1';
			M10(0) <= '1';
			M10(1) <= '1';
			--M11(0) <= '0';
			--M11(1) <= '0';
			--M12(0) <= '0';
			--M12(1) <= '0';
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '0';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0'; 
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '1' and IR(13) = '0' and IR(12) = '0') then---lw
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '1';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '1';
			M9(1) <= '1';
			M10(0) <= '0';
			M10(1) <= '0';
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= '0';
			--M12(1) <= '0';
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '0';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '0';
			Mem_en <= '1';
			Mem_R_W <= '0';
			RF_Write <= '1';
			M16(0) <= '0'; 
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
		--end if;

		elsif(IR(15) = '0' and IR(14) = '1' and IR(13) = '0' and IR(12) = '1') then---sw
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '1';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '0';
			M17 <= "00";
			M18 <= '1';
			M19 <= '1';
			M14 <= '0';
			M15 <= '0';
			Mem_en <= '1';
			Mem_R_W <= '1';
			RF_Write <= '0';
			M16(0) <= '0'; 
			M16(1) <= '0';
			M1 <= '0';
		--end if;
		
		elsif(IR(15) = '0' and IR(14) = '1' and IR(13) = '1' and IR(12) = '0') then---lm
			--M2 <= '1';
			--M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '1';
			M6 <= '1';
			M7(0) <= '0';
			M7(1) <= '1';
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(11) and IR(10) and IR(9) and M8_Control_PE;
			M10(0) <= '1';
			M10(1) <= '1';
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '0';
			Z_en <= '0';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '0';
			Mem_R_W <= '0';
			if(IR(7 downto 0) = "00000000")then
	    		Mem_en <= '0';
                        RF_Write <= '0';
	    		else
			Mem_en <= '1';
			RF_Write <= '1';
			end if;
			M16(0) <= not(addr(2) and addr(1) and addr(0)); 
			M16(1) <= '1';
			M1 <= '0';
		--end if;
		elsif(IR(15) = '0' and IR(14) = '1' and IR(13) = '1' and IR(12) = '1') then---sm
            --M2 <= '1';
            --M2 <= done;
            --PC_write_tem <= (done and HDU_output_PC);
            --IF_ID_Write <= HDU_output_IF_ID;
            --M3 <= HDU_output_M3;
	    tm20 <= '1';
            M4 <= '1';
            M5 <= '1';
            M6 <= '1';
            M7 <= "01";
            M8 <= M8_Control_PE;
            M9(0) <= '0';
            M9(1) <= IR(11) and IR(10) and IR(9) and M8_Control_PE;
            M10(0) <= '0';
            M10(1) <= addr(2) and addr(1) and addr(0);
            --M11(0) <= FDU_output;
            --M11(1) <= FDU_output;
            --M12(0) <= FDU_output;
            --M12(1) <= FDU_output;
            M13(0) <= '1';
            M13(1) <= '1';
            ALU_OP(0) <= '0';
            ALU_OP(1) <= '0';
            C_en <= '0';
            Z_en <= '0';
            M17 <= "01";
            M18 <= '1';
            M19 <= '1';
            M14 <= '1';
            M15 <= '0';
	    if(IR(7 downto 0) = "00000000")then
	    Mem_en <= '0';
            Mem_R_W <= '1';
	    else
            Mem_en <= '1';
            Mem_R_W <= '1';
	    end if;
            RF_Write <= '0';
            M16(0) <= '0'; 
            M16(1) <= '0';
            M1 <= '0';
     else
	  
	  --M2 <= done;
			--PC_write_tem <= (done and HDU_output_PC);
			--IF_ID_Write <= HDU_output_IF_ID;
			--M3 <= HDU_output_M3;
			M4 <= '0';
			M5 <= '0';
			M6 <= '0';
			M7 <= "00";
			M8 <= M8_Control_PE;
			M9(0) <= '0';
			M9(1) <= IR(5) and IR(4) and IR(3);
			M10(0) <= '0';
			M10(1) <= IR(8) and IR(7) and IR(6);
			--M11(0) <= FDU_output;
			--M11(1) <= FDU_output;
			--M12(0) <= FDU_output;
			--M12(1) <= FDU_output;
			M13(0) <= '1';
			M13(1) <= '1';
			ALU_OP(0) <= '0';
			ALU_OP(1) <= '0';
			C_en <= '1';
			Z_en <= '1';
			M17 <= "00";
			M18 <= '0';
			M19 <= '0';
			M14 <= '0';
			M15 <= '1';
			Mem_en <= '0';
			Mem_R_W <= '0';
			RF_Write <= '0';
			M16(0) <= '0';
			M16(1) <= IR(11) and IR(10) and IR(9);
			M1 <= IR(11) and IR(10) and IR(9);
	  
	  end if;
    end if;  
    end process;
PC_write <= PC_write_tem;
M2 <= M2_tem;
IF_ID_Write <= IF_ID_Write_tem;
M3 <= M3_tem;
M20 <= tm20;
end Behave;
